// bindhw5.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module bindhw5 (
		input  wire [3:0]  keys_external_connection_export, // keys_external_connection.export
		output wire [9:0]  leds_external_connection_export, // leds_external_connection.export
		input  wire        pll_ref_clk_clk,                 //              pll_ref_clk.clk
		input  wire        pll_ref_reset_reset,             //            pll_ref_reset.reset
		output wire        pll_sdram_clk_clk,               //            pll_sdram_clk.clk
		output wire [7:0]  pwm_custom_export,               //               pwm_custom.export
		output wire [12:0] sdram_wire_addr,                 //               sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                   //                         .ba
		output wire        sdram_wire_cas_n,                //                         .cas_n
		output wire        sdram_wire_cke,                  //                         .cke
		output wire        sdram_wire_cs_n,                 //                         .cs_n
		inout  wire [15:0] sdram_wire_dq,                   //                         .dq
		output wire [1:0]  sdram_wire_dqm,                  //                         .dqm
		output wire        sdram_wire_ras_n,                //                         .ras_n
		output wire        sdram_wire_we_n,                 //                         .we_n
		input  wire [9:0]  sw_external_connection_export    //   sw_external_connection.export
	);

	wire         pll_sys_clk_clk;                                             // pll:sys_clk_clk -> [KEYS:clk, LEDS:clk, SW:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_sys_clk_clk, mm_interconnect_1:pll_sys_clk_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, onchip_memory2_0:clk2, pwm_custom_0:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sysid_qsys_0:clock]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_pwm_custom_0_avalon_slave_0_chipselect;    // mm_interconnect_0:pwm_custom_0_avalon_slave_0_chipselect -> pwm_custom_0:chipselect
	wire  [31:0] mm_interconnect_0_pwm_custom_0_avalon_slave_0_readdata;      // pwm_custom_0:readdata -> mm_interconnect_0:pwm_custom_0_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_0_pwm_custom_0_avalon_slave_0_address;       // mm_interconnect_0:pwm_custom_0_avalon_slave_0_address -> pwm_custom_0:address
	wire         mm_interconnect_0_pwm_custom_0_avalon_slave_0_write;         // mm_interconnect_0:pwm_custom_0_avalon_slave_0_write -> pwm_custom_0:write
	wire  [31:0] mm_interconnect_0_pwm_custom_0_avalon_slave_0_writedata;     // mm_interconnect_0:pwm_custom_0_avalon_slave_0_writedata -> pwm_custom_0:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_keys_s1_chipselect;                        // mm_interconnect_0:KEYS_s1_chipselect -> KEYS:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                          // KEYS:readdata -> mm_interconnect_0:KEYS_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                           // mm_interconnect_0:KEYS_s1_address -> KEYS:address
	wire         mm_interconnect_0_keys_s1_write;                             // mm_interconnect_0:KEYS_s1_write -> KEYS:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                         // mm_interconnect_0:KEYS_s1_writedata -> KEYS:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                            // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                             // mm_interconnect_0:SW_s1_address -> SW:address
	wire         mm_interconnect_0_leds_s1_chipselect;                        // mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                          // LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                           // mm_interconnect_0:LEDS_s1_address -> LEDS:address
	wire         mm_interconnect_0_leds_s1_write;                             // mm_interconnect_0:LEDS_s1_write -> LEDS:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                         // mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] nios2_gen2_0_tightly_coupled_instruction_master_0_readdata;  // mm_interconnect_1:nios2_gen2_0_tightly_coupled_instruction_master_0_readdata -> nios2_gen2_0:itcm0_readdata
	wire  [27:0] nios2_gen2_0_tightly_coupled_instruction_master_0_address;   // nios2_gen2_0:itcm0_address -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_instruction_master_0_address
	wire         nios2_gen2_0_tightly_coupled_instruction_master_0_read;      // nios2_gen2_0:itcm0_read -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_instruction_master_0_read
	wire         nios2_gen2_0_tightly_coupled_instruction_master_0_clken;     // nios2_gen2_0:itcm0_clken -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_1_onchip_memory2_0_s2_chipselect;            // mm_interconnect_1:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s2_readdata;              // onchip_memory2_0:readdata2 -> mm_interconnect_1:onchip_memory2_0_s2_readdata
	wire  [15:0] mm_interconnect_1_onchip_memory2_0_s2_address;               // mm_interconnect_1:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s2_byteenable;            // mm_interconnect_1:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire         mm_interconnect_1_onchip_memory2_0_s2_write;                 // mm_interconnect_1:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s2_writedata;             // mm_interconnect_1:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_1_onchip_memory2_0_s2_clken;                 // mm_interconnect_1:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // KEYS:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [KEYS:reset_n, LEDS:reset_n, SW:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_memory2_0_reset2_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_0:reset2, pwm_custom_0:reset, rst_translator:in_reset, sdram:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         pll_reset_source_reset;                                      // pll:reset_source_reset -> rst_controller_001:reset_in0

	bindhw5_KEYS keys (
		.clk        (pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)              //                 irq.irq
	);

	bindhw5_LEDS leds (
		.clk        (pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)       // external_connection.export
	);

	bindhw5_SW sw (
		.clk      (pll_sys_clk_clk),                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_external_connection_export)     // external_connection.export
	);

	bindhw5_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_sys_clk_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	bindhw5_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_sys_clk_clk),                                            //                                  clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                                reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                                     .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //                          data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                                     .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                                     .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                                     .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                                     .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                                     .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                                     .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                                     .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //                   instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                                     .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                                     .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                                     .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                                     .readdatavalid
		.itcm0_readdata                      (nios2_gen2_0_tightly_coupled_instruction_master_0_readdata), // tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (nios2_gen2_0_tightly_coupled_instruction_master_0_address),  //                                     .address
		.itcm0_read                          (nios2_gen2_0_tightly_coupled_instruction_master_0_read),     //                                     .read
		.itcm0_clken                         (nios2_gen2_0_tightly_coupled_instruction_master_0_clken),    //                                     .clken
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                                  irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                     .writedata
		.dummy_ci_port                       ()                                                            //            custom_instruction_master.readra
	);

	bindhw5_onchip_memory2_0 onchip_memory2_0 (
		.clk         (pll_sys_clk_clk),                                  //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.address2    (mm_interconnect_1_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_1_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk2        (pll_sys_clk_clk),                                  //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                   // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	bindhw5_pll pll (
		.ref_clk_clk        (pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (pll_sdram_clk_clk),      //    sdram_clk.clk
		.reset_source_reset (pll_reset_source_reset)  // reset_source.reset
	);

	pwm pwm_custom_0 (
		.clk        (pll_sys_clk_clk),                                          //          clock.clk
		.reset      (rst_controller_reset_out_reset),                           //          reset.reset
		.address    (mm_interconnect_0_pwm_custom_0_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_pwm_custom_0_avalon_slave_0_write),      //               .write
		.chipselect (mm_interconnect_0_pwm_custom_0_avalon_slave_0_chipselect), //               .chipselect
		.writedata  (mm_interconnect_0_pwm_custom_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_pwm_custom_0_avalon_slave_0_readdata),   //               .readdata
		.pwm_out    (pwm_custom_export)                                         //        pwm_out.export
	);

	bindhw5_sdram sdram (
		.clk            (pll_sys_clk_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	bindhw5_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_sys_clk_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	bindhw5_mm_interconnect_0 mm_interconnect_0 (
		.pll_sys_clk_clk                                (pll_sys_clk_clk),                                             //                              pll_sys_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.KEYS_s1_address                                (mm_interconnect_0_keys_s1_address),                           //                                  KEYS_s1.address
		.KEYS_s1_write                                  (mm_interconnect_0_keys_s1_write),                             //                                         .write
		.KEYS_s1_readdata                               (mm_interconnect_0_keys_s1_readdata),                          //                                         .readdata
		.KEYS_s1_writedata                              (mm_interconnect_0_keys_s1_writedata),                         //                                         .writedata
		.KEYS_s1_chipselect                             (mm_interconnect_0_keys_s1_chipselect),                        //                                         .chipselect
		.LEDS_s1_address                                (mm_interconnect_0_leds_s1_address),                           //                                  LEDS_s1.address
		.LEDS_s1_write                                  (mm_interconnect_0_leds_s1_write),                             //                                         .write
		.LEDS_s1_readdata                               (mm_interconnect_0_leds_s1_readdata),                          //                                         .readdata
		.LEDS_s1_writedata                              (mm_interconnect_0_leds_s1_writedata),                         //                                         .writedata
		.LEDS_s1_chipselect                             (mm_interconnect_0_leds_s1_chipselect),                        //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.pwm_custom_0_avalon_slave_0_address            (mm_interconnect_0_pwm_custom_0_avalon_slave_0_address),       //              pwm_custom_0_avalon_slave_0.address
		.pwm_custom_0_avalon_slave_0_write              (mm_interconnect_0_pwm_custom_0_avalon_slave_0_write),         //                                         .write
		.pwm_custom_0_avalon_slave_0_readdata           (mm_interconnect_0_pwm_custom_0_avalon_slave_0_readdata),      //                                         .readdata
		.pwm_custom_0_avalon_slave_0_writedata          (mm_interconnect_0_pwm_custom_0_avalon_slave_0_writedata),     //                                         .writedata
		.pwm_custom_0_avalon_slave_0_chipselect         (mm_interconnect_0_pwm_custom_0_avalon_slave_0_chipselect),    //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.SW_s1_address                                  (mm_interconnect_0_sw_s1_address),                             //                                    SW_s1.address
		.SW_s1_readdata                                 (mm_interconnect_0_sw_s1_readdata),                            //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                         .readdata
	);

	bindhw5_mm_interconnect_1 mm_interconnect_1 (
		.pll_sys_clk_clk                                            (pll_sys_clk_clk),                                            //                                       pll_sys_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                         //          nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset2_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                             //     onchip_memory2_0_reset2_reset_bridge_in_reset.reset
		.nios2_gen2_0_tightly_coupled_instruction_master_0_address  (nios2_gen2_0_tightly_coupled_instruction_master_0_address),  // nios2_gen2_0_tightly_coupled_instruction_master_0.address
		.nios2_gen2_0_tightly_coupled_instruction_master_0_read     (nios2_gen2_0_tightly_coupled_instruction_master_0_read),     //                                                  .read
		.nios2_gen2_0_tightly_coupled_instruction_master_0_readdata (nios2_gen2_0_tightly_coupled_instruction_master_0_readdata), //                                                  .readdata
		.nios2_gen2_0_tightly_coupled_instruction_master_0_clken    (nios2_gen2_0_tightly_coupled_instruction_master_0_clken),    //                                                  .clken
		.onchip_memory2_0_s2_address                                (mm_interconnect_1_onchip_memory2_0_s2_address),              //                               onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                                  (mm_interconnect_1_onchip_memory2_0_s2_write),                //                                                  .write
		.onchip_memory2_0_s2_readdata                               (mm_interconnect_1_onchip_memory2_0_s2_readdata),             //                                                  .readdata
		.onchip_memory2_0_s2_writedata                              (mm_interconnect_1_onchip_memory2_0_s2_writedata),            //                                                  .writedata
		.onchip_memory2_0_s2_byteenable                             (mm_interconnect_1_onchip_memory2_0_s2_byteenable),           //                                                  .byteenable
		.onchip_memory2_0_s2_chipselect                             (mm_interconnect_1_onchip_memory2_0_s2_chipselect),           //                                                  .chipselect
		.onchip_memory2_0_s2_clken                                  (mm_interconnect_1_onchip_memory2_0_s2_clken)                 //                                                  .clken
	);

	bindhw5_irq_mapper irq_mapper (
		.clk           (pll_sys_clk_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (pll_sys_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (pll_reset_source_reset),                 // reset_in0.reset
		.clk            (pll_sys_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
